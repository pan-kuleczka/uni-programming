module circuit(input [3:0]i, output o);
endmodule
